module top ();
    import "DPI-C" task body();
    initial begin
        body();
    end
endmodule